erpnext.ujmd.edu.sv
uvirtualbk.ujmd.edu.sv
cdmype.ujmd.edu.sv
laboratoriosonline.ujmd.edu.sv
aulasvirtuales.ujmd.edu.sv
admisiones.ujmd.edu.sv
webquery.ujmd.edu.sv
checkout.ujmd.edu.sv
formacionc.ujmd.edu.sv
uvirtual.ujmd.edu.sv
conscius3.ujmd.edu.sv
www.conscius.ujmd.edu.sv
iij.ujmd.edu.sv
correo.ujmd.edu.sv
conscius.ujmd.edu.sv
www.ujmd.edu.sv
biblioteca.ujmd.edu.sv
itportal.ujmd.edu.sv
proyeccionsocial.ujmd.edu.sv
email.ujmd.edu.sv
beneficios.ujmd.edu.sv
conscius2.ujmd.edu.sv
medicinapaliativa.ujmd.edu.sv
cich.ujmd.edu.sv
rrhh.ujmd.edu.sv
ujmd.edu.sv
cemprende.ujmd.edu.sv
