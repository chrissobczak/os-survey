NOERROR
NOERROR
NOERROR
NOERROR
NXDOMAIN
NXDOMAIN
NOERROR
NOERROR
NOERROR
NXDOMAIN
NXDOMAIN
NXDOMAIN
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NXDOMAIN
NOERROR
NOERROR
NXDOMAIN
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NOERROR
NXDOMAIN
NXDOMAIN
NXDOMAIN
NOERROR
NOERROR
NOERROR
