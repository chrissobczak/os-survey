NA
NA
Apache
NA
LAMQ
ESF
Apache
Apache
Apache
Apache
Apache/2.4.18 (Ubuntu)
Apache
Apache
Apache
Apache/2.4.18 (Ubuntu)
Apache
Apache
ESF
Apache
ghs
ESF
Apache
ESF
Apache
Apache
Apache
Apache
